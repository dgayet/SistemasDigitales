library IEEE;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package t_types is
    type t_state is (S0, S1, S2, S3, S4, S5);
end package t_types;